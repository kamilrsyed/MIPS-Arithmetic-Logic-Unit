library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE ieee.numeric_std.ALL;


entity SYED_register_file is
port(
 rd1add			: in std_logic_vector(4 downto 0);
 rd2add			: in std_logic_vector(4 downto 0);
 wradd			: in std_logic_vector(4 downto 0);
 data				: in std_logic_vector(31 downto 0); 
 wren				: in std_logic;    
 clock			: in std_logic; 
 Q1				: out std_logic_vector(31 downto 0);
 Q2				: out std_logic_vector(31 downto 0) 
);
end SYED_register_file;

architecture Behavioral of SYED_register_file is
--initializizng memory array
type SYED_mem is array (0 to 31 ) of std_logic_vector (31 downto 0);

signal SYED_memory_array: SYED_mem:=(
	"00000000000000000100000000000000",
	"00000000000000001000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
   "00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
   "00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000", 
   "00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
   "00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
   "00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
   "00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
   "00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000"
	);

begin	
	process(clock)
	begin
	 if(rising_edge(clock)) then
	 
		 if(wren='1') then 
			--converting address to integer
		 SYED_memory_array(to_integer(unsigned(wradd))) <= data;
		 end if;
		 
	 end if;
	end process;
	
	 -- output
	 Q1 <= SYED_memory_array(to_integer(unsigned(rd1add)));
	 Q2 <= SYED_memory_array(to_integer(unsigned(rd2add)));
end Behavioral;