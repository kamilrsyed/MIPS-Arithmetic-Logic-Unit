library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE ieee.numeric_std.ALL;


entity SYED_MDR is
port(
 rdaddr			: in std_logic_vector(4 downto 0);
 wraddr			: in std_logic_vector(4 downto 0);
 data				: in std_logic_vector(31 downto 0); 
 wren				: in std_logic;    
 clock			: in std_logic; 
 Q				: out std_logic_vector(31 downto 0)
);
end SYED_MDR;

architecture Behavioral of SYED_MDR is
--initializizng memory array
type SYED_mem_MDR is array (0 to 31 ) of std_logic_vector (31 downto 0);

signal SYED_MDR_array: SYED_mem_MDR:=(
	"00000000000000000100000000000000",
	"00000000000000001000000000000000",
	"00000000000000000001110000000000",
	"00000000000000000011110000000000",
   "00000000111100000000000000000000",
	"00000000111000000100000000000000",
	"00000000000011111000000000000000",
	"00000000000000001100000000000000",
   "00000000000000111000000000000000",
	"00000000000000000000000000011000",
	"00000001110000000000000000000000",
	"00000000000000110000000000000000", 
   "00000000000000001000000000000000",
	"00000000000000000000000011100000",
	"00000000000000000000001111100000",
	"00000000000001111000000000000000",
   "00000000000000000000000000000000",
	"00000000000000000000111100001000",
	"00000011000000000000000000000000",
	"00000000000110000000000000000000",
   "00000000000000000011000000000000",
	"00000000000000001111000000000000",
	"00000000000000000000111000000000",
	"00000000000000001111000000000000",
   "00000001000000000000011000000000",
	"00000000100000001111000000000000",
	"00000010000000000000001111100000",
	"00001000000000000000000000000000",
   "00000010000000000000001111100000",
	"00100000000000000000000000000000",
	"00000100000000000000001111100000",
	"00001000000000001111000000000000"
	);

begin	
	process(clock)
	begin
	 if(rising_edge(clock)) then
	 
		 if(wren='1') then 
			--converting address to integer
		 SYED_MDR_array(to_integer(unsigned(wraddr))) <= data;
		 end if;
		 
	 end if;
	end process;
	
	 -- output
	 Q <= SYED_MDR_array(to_integer(unsigned(rdaddr)));
end Behavioral;